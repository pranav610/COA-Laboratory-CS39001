`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:35:08 10/28/2022 
// Design Name: 
// Module Name:    binary_to_bcd 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module binary_to_bcd(diff, diff_out);
	input [31:0] diff;
	output reg [5:0] diff_out;
	
	always @(*) begin
		case(diff)
			32'b10000000000000000000000000000000: diff_out = 6'd32;
			32'b01000000000000000000000000000000: diff_out = 6'd31;
			32'b00100000000000000000000000000000: diff_out = 6'd30;
			32'b00010000000000000000000000000000: diff_out = 6'd29;
			32'b00001000000000000000000000000000: diff_out = 6'd28;
			32'b00000100000000000000000000000000: diff_out = 6'd27;
			32'b00000010000000000000000000000000: diff_out = 6'd26;
			32'b00000001000000000000000000000000: diff_out = 6'd25;
			32'b00000000100000000000000000000000: diff_out = 6'd24;
			32'b00000000010000000000000000000000: diff_out = 6'd23;
			32'b00000000001000000000000000000000: diff_out = 6'd22;
			32'b00000000000100000000000000000000: diff_out = 6'd21;
			32'b00000000000010000000000000000000: diff_out = 6'd20;
			32'b00000000000001000000000000000000: diff_out = 6'd19;
			32'b00000000000000100000000000000000: diff_out = 6'd18;
			32'b00000000000000010000000000000000: diff_out = 6'd17;
			32'b00000000000000001000000000000000: diff_out = 6'd16;
			32'b00000000000000000100000000000000: diff_out = 6'd15;
			32'b00000000000000000010000000000000: diff_out = 6'd14;
			32'b00000000000000000001000000000000: diff_out = 6'd13;
			32'b00000000000000000000100000000000: diff_out = 6'd12;
			32'b00000000000000000000010000000000: diff_out = 6'd11;
			32'b00000000000000000000001000000000: diff_out = 6'd10;
			32'b00000000000000000000000100000000: diff_out = 6'd9;
			32'b00000000000000000000000010000000: diff_out = 6'd8;
			32'b00000000000000000000000001000000: diff_out = 6'd7;
			32'b00000000000000000000000000100000: diff_out = 6'd6;
			32'b00000000000000000000000000010000: diff_out = 6'd5;
			32'b00000000000000000000000000001000: diff_out = 6'd4;
			32'b00000000000000000000000000000100: diff_out = 6'd3;
			32'b00000000000000000000000000000010: diff_out = 6'd2;
			32'b00000000000000000000000000000001: diff_out = 6'd1;
			32'b00000000000000000000000000000000: diff_out = 6'd0;
			default: diff_out = 6'd0;
		endcase
	end

endmodule
