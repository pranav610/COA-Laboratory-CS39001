`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:57:31 10/19/2022 
// Design Name: 
// Module Name:    ALU 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ALU(wire a, wire b, wire less, wire Ainvert, wire Binvert, wire CarryIn, wire Operation, wire Result, wire Set, wire Overflow);
input wire a,b,less,Ainvert,Binvert,CarryIn,Operation;
output wire Result, Set, Overflow;






endmodule
